library verilog;
use verilog.vl_types.all;
entity Transmisor_vlg_check_tst is
    port(
        Salida          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Transmisor_vlg_check_tst;
