library verilog;
use verilog.vl_types.all;
entity conversor_vlg_vec_tst is
end conversor_vlg_vec_tst;
