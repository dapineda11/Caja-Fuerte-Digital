library verilog;
use verilog.vl_types.all;
entity Transmisor_vlg_vec_tst is
end Transmisor_vlg_vec_tst;
